module TotientCounter_tb

endmodule 