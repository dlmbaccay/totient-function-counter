module TotientCounter

endmodule